////////////////////////////////////////////////////////////////////////////////////////////////////////
//
// Institution   : Bandung Institute of Technology
// Engineer      : Jhonson Lee, Bobbi W. Yogatama, Hans Christian
//
// Create Date   : 11/14/2017 
// Module Name   : adder2
// Project Name  : LSI Design Contest in Okinawa 2018
// Target Devices: Sigmoid Function
// Tool versions : Vivado 2016.4
//
// Description: 
// 		Performing addition between two value
// 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: Addtion using operator +
//
///////////////////////////////////////////////////////////////////////////////////////////////////////

module adder2(a,b,c);

parameter DWIDTH=16;							
parameter AWIDTH=10;								
parameter IWIDTH=64;
parameter Layer=15;

input signed [DWIDTH-1:0] a,b;
output signed [DWIDTH-1:0] c;
assign c=a+b;
endmodule